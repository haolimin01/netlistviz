* case_1.sp simple RC 

V1 1 0 1
R1 1 2 10
R2 2 3 5
R3 3 0 1
C3 3 0 1p

.OP
.ends
