********
R1 1 0 1
R2 2 n3 2
R3 n3 0 1
IIN 1 2 1

.dc IIN 0 10 1
.end
