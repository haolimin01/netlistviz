*scale(5)	circuit type(Coupled RC tree)

VIN0 10 0 0
VIN1 11 0 1
R10 10 20 100
C10 20 0 1p
R11 11 21 100
C11 21 0 1p
*C1C 20 21 1p
R20 20 30 100
C20 30 0 1p
R21 21 31 100
C21 31 0 1p
*C2C 30 31 1p
R30 30 40 100
C30 40 0 1p
R31 31 41 100
C31 41 0 1p
*C3C 40 41 1p
R40 40 50 100
C40 50 0 1p
R41 41 51 100
C41 51 0 1p
*C4C 50 51 1p
R50 50 60 100
C50 60 0 1p
R51 51 61 100
C51 61 0 1p
*C5C 60 61 1p

.OP
.PRINT V(60) V(61)
.ENDS
