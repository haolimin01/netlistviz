* SimpleR case

V1 1 0 1
R1 1 3 1k
R2 1 2 1k
R3 2 3 1k
R4 3 0 1k
R5 2 4 1k
R6 3 5 1k
R7 0 6 1k
R8 4 5 1k
R9 5 6 1k
R10 5 7 1k
R11 4 7 1k
R12 7 6 1k
.op
.ends
